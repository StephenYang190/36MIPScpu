module Adder(x1, x2, y);
  input [29:0] x1, x2;

  output [29:0] y;

  assign y = x1 + x2;

endmodule
